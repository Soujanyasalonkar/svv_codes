module pull_try;
endmodule
