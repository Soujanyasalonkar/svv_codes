module name2;
endmodule
