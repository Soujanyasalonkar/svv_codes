module name;
endmodule
